//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : xor_gate
// File Name : xor_gate.v
// Function : Implement AND logic gate
// Designer: jessica p apuyan
// Period: Term 3 AY24-25
//-----------------------------------------------------

module xor_gate(
  input A,B,
  output C
  );
  
  // Gate type
  xor  japuyan (C, A, B);

endmodule