//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : xnor_gate
// File Name : xnor_gate.v
// Function : Implement XNOR logic gate
// Designer: Saira Cardinal
// Period: Term 3 AY24-25
//-----------------------------------------------------

module xnor_gate(
  input A,B,
  output C
  );
  
  // Gate type
  xnor scardinal (C, A, B); 

endmodule
