//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : or_gate
// File Name : or_gate.v
// Function : Implement OR logic gate
// Designer: Ernie Emago
// Period: Term 3 AY24-25
//-----------------------------------------------------

module Or_gate(
  input A,B,
  output C
  );
  
  // Gate type
  or  emago (C, A, B);

endmodule