//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : not_gate
// File Name : not_gate.v
// Function : Implement NOT logic gate
// Designer : jessica p apuyan
// Period   : Term 3 AY24-25
//-----------------------------------------------------

module not_gate(
  input A,
  output B
);

  // Gate type
  not japuyan (B, A);

endmodule