//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : xand_gate
// File Name : xand_gate.v
// Function : Implement inverse XOR (XNOR) logic gate
// Designer: Ernie Mago
// Period: Term 3 AY24-25
//-----------------------------------------------------

module xand_gate(
  input A, B,
  output C
  );

  assign C = ~(A ^ B);

endmodule
