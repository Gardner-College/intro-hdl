//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : not_gate
// File Name : not_gate.v
// Function : Implement NOT logic gate
// Designer : eric villaceran
// Period   : Term 3 AY24-25
//-----------------------------------------------------

module not_gate(
  input A,
  output B
);

  // Gate type
  not evillaceran (B, A);

endmodule
