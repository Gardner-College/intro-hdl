//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : or_gate
// File Name : or_gate.v
// Function : Implement OR logic gate
// Designer: Saira Cardinal
// Period: Term 3 AY24-25
//-----------------------------------------------------

module or_gate(
  input A,B,
  output C
  );
  
  // Gate type
  or  scardinal (C, A, B);

endmodule