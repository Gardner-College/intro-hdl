//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : xnor_gate
// File Name : xnor_gate.v
// Function : Implement AND logic gate
// Designer: Ernesto Martinez
// Period: Term 3 AY24-25
//-----------------------------------------------------

module xnor_gate(
  input A,B,
  output C
  );
  
  // Gate type
  xnor  emartinez (C, A, B);

endmodule