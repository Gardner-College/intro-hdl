//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : or_gate
// File Name : or_gate.v
// Function : Implement AND logic gate
// Designer: Ernesto T. Martinez
// Period: Term 3 AY24-25
//-----------------------------------------------------

module or_gate(
  input A,B,
  output C
  );
  
  // Gate type
  or  emartinez (C, A, B);

endmodule