//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : and_gate
// File Name : and_gate.v
// Function : Implement AND logic gate
// Designer: eric villaceran
// Period: Term 3 AY24-25
//-----------------------------------------------------

module and_gate(
  input A,B,
  output C
  );
  
  // Gate type
  and  evillaceran (C, A, B);

endmodule