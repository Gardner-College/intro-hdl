//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : xor_gate
// File Name : xor_gate.v
// Function : Implement XOR logic gate
// Designer: Ernie Mago
// Period: Term 3 AY24-25
//-----------------------------------------------------

module xor_gate(
  input A, B,
  output C
  );

  // Gate type
  xor emago (C, A, B);

endmodule
