//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name  : nor_gate
// File Name    : nor_gate.v
// Function     : Implement NOR logic gate
// Designer     : Marvin D. Llames
// Period       : Term 3 AY24-25
//-----------------------------------------------------
module nor_gate(
  input A, B,
  output C
  );

  nor MarvinL (C, A, B);

endmodule