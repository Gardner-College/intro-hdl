//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : nor_gate
// File Name : nor_gate.v
// Function : Implement AND logic gate
// Designer: Ernesto Martinez
// Period: Term 3 AY24-25
//-----------------------------------------------------

module nor_gate(
  input A,B,
  output C
  );
  
  // Gate type
  nor  emartinez (C, A, B);

endmodule