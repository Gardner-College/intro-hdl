//-----------------------------------------------------
// Laboratory Experiment 001
// Design Name : not_gate
// File Name : not_gate.v
// Function : Implement NOT logic gate
// Designer: jessica apuyan
// Period: Term 3 AY24-25
//-----------------------------------------------------

module not_gate(
  input A,
  output C
  );
  
  // Gate type
  not japuyan (C, A); 

endmodule